module TOP(port1);


	/* Island 0 */
	TSMC350nm_4x2_Indirect I__0 (.island_num(0), .row(0), .col(1), .matrix_row(1), .matrix_col(1), .Vd_P_0_row_0(net34), .Vd_P_1_row_0(net35), .Vd_P_2_row_0(net36), .Vd_P_3_row_0(net37));

 	/*Programming Mux */ 

 endmodule