VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

PROPERTYDEFINITIONS
  LAYER routingPitch REAL ;
END PROPERTYDEFINITIONS

UNITS
  DATABASE MICRONS 1000 ;
END UNITS
MANUFACTURINGGRID 0.01 ;
LAYER POLY1
  TYPE MASTERSLICE ;
END POLY1

LAYER CONT
  TYPE CUT ;
  SPACING 0.4 ;
END CONT

LAYER METAL1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0 ;
  WIDTH 0.5 ;
  SPACING 0.45 ;
  PROPERTY routingPitch 1.25 ;
END METAL1

LAYER VIA12
  TYPE CUT ;
  SPACING 0.45 ;
END VIA12

LAYER METAL2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0 ;
  WIDTH 0.6 ;
  SPACING 0.5 ;
  PROPERTY routingPitch 1.4 ;
END METAL2

LAYER VIA23
  TYPE CUT ;
  SPACING 0.45 ;
END VIA23

LAYER METAL3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0 ;
  WIDTH 0.6 ;
  SPACING 0.5 ;
  PROPERTY routingPitch 1.25 ;
END METAL3

LAYER VIA34
  TYPE CUT ;
  SPACING 0.45 ;
END VIA34

LAYER METAL4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0 ;
  WIDTH 0.6 ;
  SPACING 0.6 ;
  PROPERTY routingPitch 1.4 ;
END METAL4

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

VIARULE M4_M3 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER METAL4 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3

VIARULE M3_M2 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2

VIARULE M2_M1 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1

VIARULE M1_POLY1 GENERATE
  LAYER POLY1 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER CONT ;
    RECT -0.2 -0.2 0.2 0.2 ;
    SPACING 1 BY 1 ;
END M1_POLY1

VIA M1_POLY1
  LAYER CONT ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER POLY1 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER METAL1 ;
    RECT -0.35 -0.35 0.35 0.35 ;
END M1_POLY1

VIA M2_M1
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
  LAYER METAL2 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER METAL1 ;
    RECT -0.45 -0.45 0.45 0.45 ;
END M2_M1

VIA M3_M2
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
  LAYER METAL3 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER METAL2 ;
    RECT -0.45 -0.45 0.45 0.45 ;
END M3_M2

VIA M4_M3
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
  LAYER METAL4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER METAL3 ;
    RECT -0.45 -0.45 0.45 0.45 ;
END M4_M3


MACRO TSMC350nm_VinjDecode2to4_vtile_spacing
END TSMC350nm_VinjDecode2to4_vtile_spacing

MACRO TSMC350nm_VinjDecode2to4_vtile_D_bridge
END TSMC350nm_VinjDecode2to4_vtile_D_bridge

MACRO TSMC350nm_VinjDecode2to4_vtile
  PIN Vinj
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 7.78 11.04 9.06 11.45 ;
    END
  END Vinj
  PIN OUT<0>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 19.66 18.91 20.11 19.59 ;
    END
  END OUT<0>
  PIN OUT<1>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 19.66 13.41 20.12 14.1 ;
    END
  END OUT<1>
  PIN OUT<2>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 19.66 7.92 20.11 8.59 ;
    END
  END OUT<2>
  PIN OUT<3>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 19.66 2.41 20.11 3.09 ;
    END
  END OUT<3>
  PIN ENABLE
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 0.01 3.48 0.71 4.21 ;
    END
  END ENABLE
  PIN GND
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 19.52 5.0 20.12 5.99 ;
    END
  END GND
  PIN VINJ
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 19.15 21.56 20.05 21.96 ;
    END
  END VINJ
  PIN IN<1>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 6.56 20.89 7.5 22.0 ;
    END
  END IN<1>
  PIN IN<0>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 3.9 20.96 4.5 22.0 ;
    END
  END IN<0>
END TSMC350nm_VinjDecode2to4_vtile

MACRO TSMC350nm_VinjDecode2to4_vtile_C_bridge
END TSMC350nm_VinjDecode2to4_vtile_C_bridge

MACRO TSMC350nm_VinjDecode2to4_vtile_B_bridge
END TSMC350nm_VinjDecode2to4_vtile_B_bridge

MACRO TSMC350nm_VinjDecode2to4_vtile_A_bridge
END TSMC350nm_VinjDecode2to4_vtile_A_bridge

MACRO TSMC350nm_drainSelect_progrundrains
  PIN prog_drain<3>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 30.93 0.93 31.86 1.43 ;
    END
  END prog_drain<3>
  PIN prog_drain<2>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 30.97 9.62 31.86 10.12 ;
    END
  END prog_drain<2>
  PIN prog_drain<1>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 31.0 13.97 31.86 14.47 ;
    END
  END prog_drain<1>
  PIN run_drain<3>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 31.01 2.45 31.86 2.95 ;
    END
  END run_drain<3>
  PIN run_drain<2>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 30.94 5.31 31.86 5.81 ;
    END
  END run_drain<2>
  PIN prog_drain<0>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 31.12 20.75 31.86 21.25 ;
    END
  END prog_drain<0>
  PIN GND
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 4.19 21.33 4.99 22.0 ;
    END
  END GND
  PIN VINJ
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 1.4 21.5 2.8 22.0 ;
    END
  END VINJ
  PIN run_drain<0>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 31.01 19.56 31.86 20.06 ;
    END
  END run_drain<0>
  PIN run_drain<1>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 31.04 16.75 31.86 17.24 ;
    END
  END run_drain<1>
  PIN SELECT<3>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 0.0 2.54 0.67 2.97 ;
    END
  END SELECT<3>
  PIN SELET<2>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 0.0 8.03 0.67 8.46 ;
    END
  END SELET<2>
  PIN SELECT<1>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 0.0 13.54 0.67 13.97 ;
    END
  END SELECT<1>
  PIN SELECT<0>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 0.0 18.9 0.67 19.6 ;
    END
  END SELECT<0>
  PIN VINJ_b
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 21.94 0.0 23.29 0.58 ;
    END
  END VINJ_b
  PIN GND_b
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 17.16 0.0 18.16 0.58 ;
    END
  END GND_b
  PIN run_drainrail
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 27.01 21.19 27.71 22.0 ;
    END
  END run_drainrail
  PIN prog_drainrail
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 7.36 21.34 8.16 22.0 ;
    END
  END prog_drainrail
END TSMC350nm_drainSelect_progrundrains

MACRO TSMC350nm_4TGate_ST_draincutoff
  PIN In<0>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 9.96 17.5 10.6 18.45 ;
    END
  END In<0>
  PIN In<1>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 9.91 14.7 10.6 15.93 ;
    END
  END In<1>
  PIN In<2>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 10.01 6.9 10.6 7.8 ;
    END
  END In<2>
  PIN In<3>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 10.02 3.5 10.6 4.3 ;
    END
  END In<3>
  PIN A<0>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 0.0 19.56 1.4 20.06 ;
    END
  END A<0>
  PIN A<1>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 0.0 16.75 1.4 17.25 ;
    END
  END A<1>
  PIN A<2>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 0.0 5.3 1.4 5.8 ;
    END
  END A<2>
  PIN A<3>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 0.0 2.45 1.4 2.95 ;
    END
  END A<3>
  PIN P<0>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 0.0 20.75 1.4 21.25 ;
    END
  END P<0>
  PIN P<1>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 0.0 13.97 1.4 14.47 ;
    END
  END P<1>
  PIN P<2>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 0.0 9.62 1.4 10.12 ;
    END
  END P<2>
  PIN P<3>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 0.0 0.93 1.4 1.43 ;
    END
  END P<3>
  PIN PR<0>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 10.0 20.3 10.6 21.25 ;
    END
  END PR<0>
  PIN PR<1>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 10.13 11.9 10.6 12.8 ;
    END
  END PR<1>
  PIN PR<2>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 10.0 9.4 10.6 10.3 ;
    END
  END PR<2>
  PIN PR<3>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 10.0 0.7 10.6 1.6 ;
    END
  END PR<3>
  PIN VDD_b
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 7.89 0.0 8.79 0.54 ;
    END
  END VDD_b
  PIN RUN
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 5.9 21.13 6.5 22.0 ;
    END
  END RUN
  PIN VDD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 7.89 21.3 8.79 22.0 ;
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 3.35 21.3 4.25 22.0 ;
    END
  END GND
  PIN GND_b
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 3.35 0.0 4.25 0.73 ;
    END
  END GND_b
  PIN RUN_b
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 5.9 0.0 6.5 0.71 ;
    END
  END RUN_b
END TSMC350nm_4TGate_ST_draincutoff

MACRO TSMC350nm_Amplifier9T_FGBias
  PIN VD_P
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 0.0 16.87 1.4 18.27 ;
    END
  END VD_P
  PIN Vout
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 58.96 1.09 60.36 2.49 ;
    END
  END Vout
  PIN VIN_PLUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 0.0 2.76 1.4 4.16 ;
    END
  END VIN_PLUS
  PIN VD_R
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 0.0 11.17 1.4 12.57 ;
    END
  END VD_R
  PIN VIN_MINUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 0.0 6.97 1.4 8.37 ;
    END
  END VIN_MINUS
  PIN GND_b
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 51.59 0.0 52.99 1.4 ;
    END
  END GND_b
  PIN VPWR
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 42.13 20.61 43.53 22.0 ;
    END
  END VPWR
  PIN Vsel_b
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 0.66 0.0 2.06 1.4 ;
    END
  END Vsel_b
  PIN VINJ_b
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 13.85 0.0 15.25 1.4 ;
    END
  END VINJ_b
  PIN Vg_b
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 9.06 0.0 10.46 1.4 ;
    END
  END Vg_b
  PIN PROG_b
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 6.26 0.0 7.66 1.4 ;
    END
  END PROG_b
  PIN VTUN_b
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 3.46 0.0 4.86 1.4 ;
    END
  END VTUN_b
  PIN PROG
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 6.26 20.6 7.66 22.0 ;
    END
  END PROG
  PIN VINJ
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 13.85 20.6 15.25 22.0 ;
    END
  END VINJ
  PIN Vg
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 9.06 20.6 10.46 22.0 ;
    END
  END Vg
  PIN VTUN
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 3.46 20.6 4.86 22.0 ;
    END
  END VTUN
  PIN Vsel
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 0.66 20.6 2.06 22.0 ;
    END
  END Vsel
  PIN GND
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 51.59 20.6 52.99 22.0 ;
    END
  END GND
  PIN VPWR_b
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 42.13 0.01 43.53 1.4 ;
    END
  END VPWR_b
END TSMC350nm_Amplifier9T_FGBias

MACRO TSMC350nm_IndirectSwitches
  PIN GND_T
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 15.4 21.0 16.2 22.0 ;
    END
  END GND_T
  PIN VINJ_T
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 6.3 21.04 7.32 22.0 ;
    END
  END VINJ_T
  PIN VDD<1>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 24.5 0.0 25.1 0.75 ;
    END
  END VDD<1>
  PIN VTUN
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 13.3 0.0 13.9 0.82 ;
    END
  END VTUN
  PIN GND<0>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 11.2 0.0 11.8 0.85 ;
    END
  END GND<0>
  PIN GNDV<1>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 15.47 0.0 15.95 1.0 ;
    END
  END GNDV<1>
  PIN VINJ
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 4.2 0.0 4.8 1.0 ;
    END
  END VINJ
  PIN VDD<0>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 2.1 0.0 2.7 1.09 ;
    END
  END VDD<0>
  PIN Vg<0>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 8.4 0.005 9.0 0.825 ;
    END
  END Vg<0>
  PIN CTRL_B<0>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 6.3 0.01 6.9 0.76 ;
    END
  END CTRL_B<0>
  PIN CTRL_B<1>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 20.3 0.01 20.9 0.75 ;
    END
  END CTRL_B<1>
  PIN Vg<1>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 18.2 0.0 18.8 0.76 ;
    END
  END Vg<1>
  PIN decode<0>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 3.46 21.16 4.8 22.0 ;
    END
  END decode<0>
  PIN RUN_IN<1>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 17.5 21.01 18.1 22.0 ;
    END
  END RUN_IN<1>
  PIN RUN_IN<0>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 10.5 20.9 11.1 22.0 ;
    END
  END RUN_IN<0>
  PIN VPWR<1>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 21.7 21.08 22.3 22.0 ;
    END
  END VPWR<1>
  PIN decode<1>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 23.8 21.09 25.0 22.0 ;
    END
  END decode<1>
  PIN VPWR<0>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 1.71 21.21 2.43 22.0 ;
    END
  END VPWR<0>
  PIN VTUN_T
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 12.6 21.12 13.7 22.0 ;
    END
  END VTUN_T
  PIN vtun_l
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 0.0 0.9 1.31 1.88 ;
    END
  END vtun_l
  PIN vtun_r
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 26.17 0.9 27.46 2.17 ;
    END
  END vtun_r
  PIN vgsel_r
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 26.52 3.15 27.46 4.45 ;
    END
  END vgsel_r
  PIN prog_r
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 26.59 9.15 27.46 10.55 ;
    END
  END prog_r
  PIN run_r
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 26.28 6.05 27.46 7.29 ;
    END
  END run_r
  PIN RUN
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 0.0 6.05 0.91 7.29 ;
    END
  END RUN
  PIN PROG
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 0.0 9.15 0.87 10.55 ;
    END
  END PROG
  PIN Vgsel
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 0.0 3.72 0.91 4.45 ;
    END
  END Vgsel
END TSMC350nm_IndirectSwitches

MACRO TSMC350nm_VinjDecode2to4_htile
  PIN IN<1>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 0.0 11.85 0.9 12.74 ;
    END
  END IN<1>
  PIN IN<0>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 0.0 10.13 0.87 11.1 ;
    END
  END IN<0>
  PIN VINJ
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 0.0 1.99 0.5 2.49 ;
    END
  END VINJ
  PIN GND
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 0.0 6.99 0.51 7.49 ;
    END
  END GND
  PIN GND_b<1>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 40.32 0.0 40.92 1.79 ;
    END
  END GND_b<1>
  PIN VINJ_b<1>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 22.1 0.0 22.7 1.44 ;
    END
  END VINJ_b<1>
  PIN GND_b<0>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 18.85 0.0 19.45 1.41 ;
    END
  END GND_b<0>
  PIN VINJ_b<0>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 1.07 0.0 1.67 1.25 ;
    END
  END VINJ_b<0>
  PIN VINJV
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 23.7 21.26 24.31 22.0 ;
    END
  END VINJV
  PIN GNDV
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 25.84 21.28 26.44 22.0 ;
    END
  END GNDV
  PIN RUN_OUT<3>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 34.39 0.0 35.19 0.86 ;
    END
  END RUN_OUT<3>
  PIN RUN_OUT<2>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 28.77 0.0 29.57 0.86 ;
    END
  END RUN_OUT<2>
  PIN RUN_OUT<1>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 13.5 0.0 14.1 0.86 ;
    END
  END RUN_OUT<1>
  PIN RUN_OUT<0>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 7.34 0.0 8.14 0.86 ;
    END
  END RUN_OUT<0>
  PIN ENABLE
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 6.29 21.66 6.89 22.0 ;
    END
  END ENABLE
  PIN OUT<2>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 25.28 0.0 25.87 0.87 ;
    END
  END OUT<2>
  PIN OUT<3>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 37.14 0.0 37.73 0.83 ;
    END
  END OUT<3>
  PIN OUT<0>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 4.27 0.0 4.87 0.86 ;
    END
  END OUT<0>
  PIN OUT<1>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 16.14 0.0 16.72 0.85 ;
    END
  END OUT<1>
  PIN VGRUN<0>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 9.1 21.59 9.7 22.0 ;
    END
  END VGRUN<0>
  PIN VGRUN<1>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 11.2 21.6 11.8 22.0 ;
    END
  END VGRUN<1>
  PIN VGRUN<2>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 28.7 21.71 29.3 22.0 ;
    END
  END VGRUN<2>
  PIN VGRUN<3>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 33.6 21.54 34.2 22.0 ;
    END
  END VGRUN<3>
END TSMC350nm_VinjDecode2to4_htile

MACRO TGate_DT
  PIN SELA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 0.0 13.5 1.4 14.9 ;
    END
  END SELA
  PIN C
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 0.0 6.78 1.4 8.18 ;
    END
  END C
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 7.18 9.11 8.58 10.51 ;
    END
  END B
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 7.18 14.37 8.58 15.77 ;
    END
  END A
  PIN VDD_b
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 4.07 0.0 5.47 1.4 ;
    END
  END VDD_b
  PIN GND_b
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 1.82 0.0 3.22 1.4 ;
    END
  END GND_b
  PIN GND
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 1.82 20.6 3.22 22.0 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 4.07 20.6 5.47 22.0 ;
    END
  END VDD
END TGate_DT

MACRO Capacitor_80ff
  PIN Bot
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 20.21 10.47 21.31 12.17 ;
    END
  END Bot
  PIN Top
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 0.0 10.48 1.16 12.17 ;
    END
  END Top
END Capacitor_80ff

MACRO tile_analog_frame
  PIN n_Prog
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 13.3 285.6 14.7 288.4 ;
    END
  END n_Prog
  PIN n_Run
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 27.3 285.6 28.7 288.4 ;
    END
  END n_Run
  PIN n_AVDD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 41.3 285.6 42.7 288.4 ;
    END
  END n_AVDD
  PIN n_gnd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 313.91 285.6 315.31 288.4 ;
    END
  END n_gnd
  PIN n_vinj
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 299.91 285.6 301.31 288.4 ;
    END
  END n_vinj
  PIN n_RST
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 55.3 285.6 56.7 288.4 ;
    END
  END n_RST
  PIN n_Code<0>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 69.3 285.6 70.7 288.4 ;
    END
  END n_Code<0>
  PIN n_Code<1>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 83.3 285.6 84.7 288.4 ;
    END
  END n_Code<1>
  PIN n_Code<2>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 97.3 285.6 98.7 288.4 ;
    END
  END n_Code<2>
  PIN n_Code<3>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 111.3 285.6 112.7 288.4 ;
    END
  END n_Code<3>
  PIN n_Code<4>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 125.3 285.6 126.7 288.4 ;
    END
  END n_Code<4>
  PIN s_gnd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 313.91 0.0 315.31 2.8 ;
    END
  END s_gnd
  PIN s_vinj
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 299.91 0.0 301.31 2.8 ;
    END
  END s_vinj
  PIN s_Vout
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 13.3 0.0 14.7 2.8 ;
    END
  END s_Vout
  PIN w_DrainB<0>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 273.0 2.8 274.4 ;
    END
  END w_DrainB<0>
  PIN w_DrainB<1>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 259.0 2.8 260.4 ;
    END
  END w_DrainB<1>
  PIN w_DrainB<2>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 245.0 2.8 246.4 ;
    END
  END w_DrainB<2>
  PIN w_DrainB<3>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 231.0 2.8 232.4 ;
    END
  END w_DrainB<3>
  PIN w_DrainEnable
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 217.0 2.8 218.4 ;
    END
  END w_DrainEnable
  PIN w_GateB<0>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 203.0 2.8 204.4 ;
    END
  END w_GateB<0>
  PIN w_GateB<1>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 189.0 2.8 190.4 ;
    END
  END w_GateB<1>
  PIN w_GateEnable
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 0.0 175.0 2.8 176.4 ;
    END
  END w_GateEnable
END tile_analog_frame

MACRO EPOT
  PIN Vout
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 83.26 0.74 84.76 2.14 ;
    END
  END Vout
  PIN Vd_P<1>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 0.0 2.09 1.4 3.39 ;
    END
  END Vd_P<1>
  PIN Vd_P<0>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 0.0 18.35 1.4 19.65 ;
    END
  END Vd_P<0>
  PIN Vin+
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 0.0 13.78 1.4 15.08 ;
    END
  END Vin+
  PIN GND_b
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 76.77 0.0 78.17 1.4 ;
    END
  END GND_b
  PIN VDD_b
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 39.68 0.0 41.08 1.4 ;
    END
  END VDD_b
  PIN Vg_b<1>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 35.5 0.0 36.9 1.4 ;
    END
  END Vg_b<1>
  PIN Vsel_b<1>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 28.93 0.0 30.33 1.4 ;
    END
  END Vsel_b<1>
  PIN Prog_b
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 26.08 0.0 27.48 1.4 ;
    END
  END Prog_b
  PIN VTUN_b
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 21.4 0.0 22.8 1.4 ;
    END
  END VTUN_b
  PIN Vg_b<0>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 18.37 0.0 19.77 1.4 ;
    END
  END Vg_b<0>
  PIN Vsel_b<0>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 3.6 0.0 5.0 1.4 ;
    END
  END Vsel_b<0>
  PIN VINJ_b
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 1.04 0.0 2.44 1.4 ;
    END
  END VINJ_b
  PIN Vg<1>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 35.5 20.6 36.9 22.0 ;
    END
  END Vg<1>
  PIN VTUN
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 21.4 20.6 22.8 22.0 ;
    END
  END VTUN
  PIN Vsel<0>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 3.6 20.6 5.0 22.0 ;
    END
  END Vsel<0>
  PIN GND
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 76.77 20.6 78.17 22.0 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 39.68 20.6 41.08 22.0 ;
    END
  END VDD
  PIN Prog
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 26.08 20.6 27.48 22.0 ;
    END
  END Prog
  PIN Vg<0>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 18.37 20.6 19.77 22.0 ;
    END
  END Vg<0>
  PIN VINJ
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 1.04 20.6 2.44 22.0 ;
    END
  END VINJ
  PIN Vsel<1>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 28.93 20.6 30.33 22.0 ;
    END
  END Vsel<1>
END EPOT

END LIBRARY