module TOP(port1);


	/* Island 0 */
	TSMC350nm_TA2Cell_Weak I__0 (.island_num(0), .row(0), .col(0), .matrix_row(1), .matrix_col(1), .VD_P_0_row_0(net222[0]), .VD_P_1_row_0(net223[0]), .VIN1_PLUSrow_0(net298), .VIN1_MINUSrow_0(net30), .VIN2_PLUSrow_0(net30), .VIN2_MINUSrow_0(net71), .OUTPUT_0_row_0(net30), .OUTPUT_1_row_0(net30), .Vsel_0_row_0(net296), .Vsel_1_row_0(net297), .RUNrow_0(net325), .Vg_0_row_0(net294), .Vg_1_row_0(net295), .PROGrow_0(net324), .VTUNrow_0(net322), .VINJrow_0(net320), .GNDrow_0(net321), .VPWRrow_0(net323));
	TSMC350nm_TA2Cell_Weak I__1 (.island_num(0), .row(1), .col(0), .matrix_row(1), .matrix_col(1), .VD_P_0_row_0(net224[0]), .VD_P_1_row_0(net225[0]), .VIN1_PLUSrow_0(net30), .VIN1_MINUSrow_0(net71), .VIN2_PLUSrow_0(net71), .VIN2_MINUSrow_0(net300), .OUTPUT_0_row_0(net71), .OUTPUT_1_row_0(net300));
	TSMC350nm_TA2Cell_Weak I__2 (.island_num(0), .row(2), .col(0), .matrix_row(1), .matrix_col(1), .VD_P_0_row_0(net226[0]), .VD_P_1_row_0(net227[0]), .VIN1_PLUSrow_0(net71), .VIN1_MINUSrow_0(net72), .VIN2_PLUSrow_0(net72), .VIN2_MINUSrow_0(net113), .OUTPUT_0_row_0(net72), .OUTPUT_1_row_0(net72));
	TSMC350nm_TA2Cell_Weak I__3 (.island_num(0), .row(3), .col(0), .matrix_row(1), .matrix_col(1), .VD_P_0_row_0(net228[0]), .VD_P_1_row_0(net229[0]), .VIN1_PLUSrow_0(net72), .VIN1_MINUSrow_0(net113), .VIN2_PLUSrow_0(net113), .VIN2_MINUSrow_0(net301), .OUTPUT_0_row_0(net113), .OUTPUT_1_row_0(net301));
	TSMC350nm_TA2Cell_Weak I__4 (.island_num(0), .row(4), .col(0), .matrix_row(1), .matrix_col(1), .VD_P_0_row_0(net230[0]), .VD_P_1_row_0(net231[0]), .VIN1_PLUSrow_0(net113), .VIN1_MINUSrow_0(net114), .VIN2_PLUSrow_0(net114), .VIN2_MINUSrow_0(net155), .OUTPUT_0_row_0(net114), .OUTPUT_1_row_0(net114));
	TSMC350nm_TA2Cell_Weak I__5 (.island_num(0), .row(5), .col(0), .matrix_row(1), .matrix_col(1), .VD_P_0_row_0(net232[0]), .VD_P_1_row_0(net233[0]), .VIN1_PLUSrow_0(net114), .VIN1_MINUSrow_0(net155), .VIN2_PLUSrow_0(net155), .VIN2_MINUSrow_0(net302), .OUTPUT_0_row_0(net155), .OUTPUT_1_row_0(net302));
	TSMC350nm_TA2Cell_Weak I__6 (.island_num(0), .row(6), .col(0), .matrix_row(1), .matrix_col(1), .VD_P_0_row_0(net234[0]), .VD_P_1_row_0(net235[0]), .VIN1_PLUSrow_0(net155), .VIN1_MINUSrow_0(net156), .VIN2_PLUSrow_0(net156), .VIN2_MINUSrow_0(net195), .OUTPUT_0_row_0(net156), .OUTPUT_1_row_0(net156));
	TSMC350nm_TA2Cell_Weak I__7 (.island_num(0), .row(7), .col(0), .matrix_row(1), .matrix_col(1), .VD_P_0_row_0(net236[0]), .VD_P_1_row_0(net237[0]), .VIN1_PLUSrow_0(net156), .VIN1_MINUSrow_0(net195), .VIN2_PLUSrow_0(net195), .VIN2_MINUSrow_0(net303), .OUTPUT_0_row_0(net195), .OUTPUT_1_row_0(net303));
	TSMC350nm_TA2Cell_Weak I__8 (.island_num(0), .row(8), .col(0), .matrix_row(1), .matrix_col(1), .VD_P_0_row_0(net238[0]), .VD_P_1_row_0(net239[0]), .VIN1_PLUSrow_0(net195), .VIN1_MINUSrow_0(net196), .VIN2_PLUSrow_0(net196), .VIN2_MINUSrow_0(net299), .OUTPUT_0_row_0(net196), .OUTPUT_1_row_0(net196));
	TSMC350nm_TA2Cell_Weak I__9 (.island_num(0), .row(9), .col(0), .matrix_row(1), .matrix_col(1), .VD_P_0_row_0(net240[0]), .VD_P_1_row_0(net241[0]), .VIN1_PLUSrow_0(net196), .VIN1_MINUSrow_0(net299), .VIN2_PLUSrow_0(net299), .VIN2_MINUSrow_0(net304), .OUTPUT_0_row_0(net299), .OUTPUT_1_row_0(net304), .VINJ_brow_0(net319), .GND_brow_0(net318));

 	/*Programming Mux */ 
	TSMC350nm_VinjDecode2to4_vtile decoder(.island_num(0), .direction(vertical), .bits(5), .decode_n0_VINJ(net319), .decode_n0_GND(net318), .decode_n0_IN_0_(net316), .decode_n2_IN_1_(net315), .decode_n2_IN_0_(net314), .decode_n4_IN_1_(net313), .decode_n4_IN_0_(net312), .decode_n0_ENABLE(net317));
	TSMC350nm_drainSelect_progrundrains switch(.island_num(0), .direction(vertical), .num(5), .type(drain_select), .switch_n0_prog_drainrail(net311), .switch_n0_VINJ(net319), .switch_n0_GND(net318));
	TSMC350nm_4TGate_ST_draincutoff switch(.island_num(0), .direction(vertical), .num(5), .type(prog_switch), .switch_n0_PR_0_(net222[0]), .switch_n0_PR_1_(net223[0]), .switch_n0_PR_2_(net224[0]), .switch_n0_PR_3_(net225[0]), .switch_n1_PR_0_(net226[0]), .switch_n1_PR_1_(net227[0]), .switch_n1_PR_2_(net228[0]), .switch_n1_PR_3_(net229[0]), .switch_n2_PR_0_(net230[0]), .switch_n2_PR_1_(net231[0]), .switch_n2_PR_2_(net232[0]), .switch_n2_PR_3_(net233[0]), .switch_n3_PR_0_(net234[0]), .switch_n3_PR_1_(net235[0]), .switch_n3_PR_2_(net236[0]), .switch_n3_PR_3_(net237[0]), .switch_n4_PR_0_(net238[0]), .switch_n4_PR_1_(net239[0]), .switch_n4_PR_2_(net240[0]), .switch_n4_PR_3_(net241[0]), .switch_n0_VDD(net319), .switch_n0_GND(net318), .switch_n0_RUN(net325));
	TSMC350nm_VinjDecode2to4_htile decoder(.island_num(0), .direction(horizontal), .bits(2), .decode_n0_ENABLE(net308), .decode_n0_VINJ_b_0_(net306), .decode_n0_VINJV(net320), .decode_n0_GNDV(net321), .decode_n0_n0_IN_1_(net310), .decode_n0_n0_IN_0_(net309));
	TSMC350nm_IndirectSwitches switch(.island_num(0), .direction(horizontal), .num(1), .switch_n0_GND_T(net321), .switch_n0_VINJ_T(net306), .switch_n0_CTRL_B_0_(net296), .switch_n0_CTRL_B_1_(net297), .switch_n0_Vg_0_(net294), .switch_n0_Vg_1_(net295));
	TSMC350nm_IndirectSwitches switch_ind(.island_num(0), .direction(horizontal), .col(0), .RUN_IN_0_(net305), .RUN_IN_1_(net305), .PROG(net324), .RUN(net325), .Vgsel(net307));


	/* Frame */ 
	tile_analog_frame cab_frame(.pin_layer(METAL3), .W_w_Vin(net298), .E_e_Vout(net299), .E_e_Vout_Buf_0_(net300), .E_e_Vout_Buf_1_(net301), .E_e_Vout_Buf_2_(net302), .E_e_Vout_Buf_3_(net303), .E_e_Vout_Buf_4_(net304), .N_n_Prog(net324), .N_n_Run(net325), .N_n_VGRUN(net305), .N_n_VGPROG(net307), .N_n_VTUN(net322), .N_n_AVDD(net323), .N_n_gnd(net321), .S_s_gnd(net318), .N_n_vinj(net320), .S_s_vinj(net319), .S_s_Drainline_Prog(net311), .N_n_GateEnable(net308), .W_w_GateB_0_(net309), .W_w_GateB_1_(net310), .W_w_DrainEnable(net317), .W_w_DrainB_0_(net312), .W_w_DrainB_1_(net313), .W_w_DrainB_2_(net314), .W_w_DrainB_3_(net315), .W_w_DrainB_4_(net316));
 endmodule