VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

PROPERTYDEFINITIONS
  LAYER routingPitch REAL ;
END PROPERTYDEFINITIONS

UNITS
  DATABASE MICRONS 1000 ;
END UNITS
MANUFACTURINGGRID 0.01 ;
LAYER POLY1
  TYPE MASTERSLICE ;
END POLY1

LAYER CONT
  TYPE CUT ;
  SPACING 0.4 ;
END CONT

LAYER METAL1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0 ;
  WIDTH 0.5 ;
  SPACING 0.45 ;
  PROPERTY routingPitch 1.25 ;
END METAL1

LAYER VIA12
  TYPE CUT ;
  SPACING 0.45 ;
END VIA12

LAYER METAL2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0 ;
  WIDTH 0.6 ;
  SPACING 0.5 ;
  PROPERTY routingPitch 1.4 ;
END METAL2

LAYER VIA23
  TYPE CUT ;
  SPACING 0.45 ;
END VIA23

LAYER METAL3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0 ;
  WIDTH 0.6 ;
  SPACING 0.5 ;
  PROPERTY routingPitch 1.25 ;
END METAL3

LAYER VIA34
  TYPE CUT ;
  SPACING 0.45 ;
END VIA34

LAYER METAL4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0 ;
  WIDTH 0.6 ;
  SPACING 0.6 ;
  PROPERTY routingPitch 1.4 ;
END METAL4

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

VIARULE M4_M3 GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER METAL4 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M4_M3

VIARULE M3_M2 GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER METAL3 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M3_M2

VIARULE M2_M1 GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER METAL2 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1 BY 1 ;
END M2_M1

VIARULE M1_POLY1 GENERATE
  LAYER POLY1 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER METAL1 ;
    ENCLOSURE 0.15 0.15 ;
  LAYER CONT ;
    RECT -0.2 -0.2 0.2 0.2 ;
    SPACING 1 BY 1 ;
END M1_POLY1

VIA M1_POLY1
  LAYER CONT ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER POLY1 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER METAL1 ;
    RECT -0.35 -0.35 0.35 0.35 ;
END M1_POLY1

VIA M2_M1
  LAYER VIA12 ;
    RECT -0.25 -0.25 0.25 0.25 ;
  LAYER METAL2 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER METAL1 ;
    RECT -0.45 -0.45 0.45 0.45 ;
END M2_M1

VIA M3_M2
  LAYER VIA23 ;
    RECT -0.25 -0.25 0.25 0.25 ;
  LAYER METAL3 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER METAL2 ;
    RECT -0.45 -0.45 0.45 0.45 ;
END M3_M2

VIA M4_M3
  LAYER VIA34 ;
    RECT -0.25 -0.25 0.25 0.25 ;
  LAYER METAL4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER METAL3 ;
    RECT -0.45 -0.45 0.45 0.45 ;
END M4_M3


MACRO TSMC350nm_4x2_Indirect
  PIN Vg<1>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 18.2 21.06 18.8 22.0 ;
    END
  END Vg<1>
  PIN Vsel<1>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 20.3 21.08 20.9 22.0 ;
    END
  END Vsel<1>
  PIN VINJ<1>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 22.4 21.05 23.0 22.0 ;
    END
  END VINJ<1>
  PIN Vsel<0>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 6.3 21.2 6.9 22.0 ;
    END
  END Vsel<0>
  PIN Vs<0>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 2.1 21.21 2.7 22.0 ;
    END
  END Vs<0>
  PIN Vs<1>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 24.5 21.06 25.1 22.0 ;
    END
  END Vs<1>
  PIN VTUN
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 13.3 21.09 13.9 22.0 ;
    END
  END VTUN
  PIN VINJ<0>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 4.2 21.18 4.8 22.0 ;
    END
  END VINJ<0>
  PIN GND<0>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 11.2 21.07 11.8 22.0 ;
    END
  END GND<0>
  PIN Vg<0>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 8.4 21.03 9.0 22.0 ;
    END
  END Vg<0>
  PIN GND<1>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 15.41 21.06 16.01 22.0 ;
    END
  END GND<1>
  PIN Vs_b<0>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 1.42 0.0 2.7 0.6 ;
    END
  END Vs_b<0>
  PIN VINJ_b<0>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 4.2 0.0 4.8 0.76 ;
    END
  END VINJ_b<0>
  PIN Vsel_b<0>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 6.3 0.0 6.9 0.78 ;
    END
  END Vsel_b<0>
  PIN Vg_b<0>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 8.4 0.0 9.0 0.77 ;
    END
  END Vg_b<0>
  PIN GND_b<0>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 11.2 0.0 11.8 0.76 ;
    END
  END GND_b<0>
  PIN VTUN_b
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 13.3 0.0 13.9 0.76 ;
    END
  END VTUN_b
  PIN GND_b<1>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 15.41 0.0 16.01 0.83 ;
    END
  END GND_b<1>
  PIN Vg_b<1>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 18.2 0.0 18.8 0.76 ;
    END
  END Vg_b<1>
  PIN Vsel_b<1>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 20.3 0.0 20.9 0.75 ;
    END
  END Vsel_b<1>
  PIN VINJ_b<1>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 22.4 0.0 23.0 0.77 ;
    END
  END VINJ_b<1>
  PIN Vs_b<1>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 24.5 0.0 25.75 0.61 ;
    END
  END Vs_b<1>
  PIN Vd_Pl<3>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 0.0 0.7 1.47 1.2 ;
    END
  END Vd_Pl<3>
  PIN Vd_Rl<3>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 0.0 3.5 1.45 4.0 ;
    END
  END Vd_Rl<3>
  PIN Vd_Rl<2>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 0.0 7.0 1.4 7.5 ;
    END
  END Vd_Rl<2>
  PIN Vd_Pl<2>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 0.0 9.8 1.41 10.3 ;
    END
  END Vd_Pl<2>
  PIN Vd_Pl<1>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 0.0 11.89 1.43 12.4 ;
    END
  END Vd_Pl<1>
  PIN Vd_Rl<1>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 0.0 14.7 1.46 15.2 ;
    END
  END Vd_Rl<1>
  PIN Vd_Rl<0>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 0.0 17.5 1.43 18.0 ;
    END
  END Vd_Rl<0>
  PIN Vd_Pl<0>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 0.0 20.3 1.4 20.9 ;
    END
  END Vd_Pl<0>
  PIN Vd_P<0>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 26.63 20.3 27.46 20.8 ;
    END
  END Vd_P<0>
  PIN Vd_R<1>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 26.56 14.7 27.44 15.2 ;
    END
  END Vd_R<1>
  PIN Vd_R<3>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 26.5 3.5 27.46 4.0 ;
    END
  END Vd_R<3>
  PIN Vd_P<3>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 26.55 0.7 27.46 1.2 ;
    END
  END Vd_P<3>
  PIN Vd_P<1>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 26.38 11.9 27.46 12.4 ;
    END
  END Vd_P<1>
  PIN Vd_P<2>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 26.51 9.8 27.46 10.3 ;
    END
  END Vd_P<2>
  PIN Vd_R<0>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 26.66 17.5 27.46 18.0 ;
    END
  END Vd_R<0>
  PIN Vd_R<2>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 26.53 7.0 27.46 7.5 ;
    END
  END Vd_R<2>
END TSMC350nm_4x2_Indirect

MACRO dotproduct_R
  PIN GND
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 14.71 21.4 15.31 22.0 ;
    END
  END GND
  PIN out2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 17.05 21.4 17.65 22.0 ;
    END
  END out2
  PIN out1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 6.95 21.4 7.55 22.0 ;
    END
  END out1
  PIN phi2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 11.45 21.4 12.05 22.0 ;
    END
  END phi2
  PIN phi1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 2.1 21.4 2.7 22.0 ;
    END
  END phi1
  PIN Q<0>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 0.0 16.61 1.4 18.01 ;
    END
  END Q<0>
  PIN Q<3>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 0.0 4.01 1.4 5.41 ;
    END
  END Q<3>
  PIN Q<1>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 0.0 14.76 1.4 16.16 ;
    END
  END Q<1>
  PIN Q<2>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 0.0 5.86 1.4 7.26 ;
    END
  END Q<2>
  PIN K<2>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 20.6 7.01 22.0 8.41 ;
    END
  END K<2>
  PIN K<1>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 20.6 13.81 22.0 15.21 ;
    END
  END K<1>
  PIN K<3>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 20.6 2.61 22.0 4.01 ;
    END
  END K<3>
  PIN K<0>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 20.6 17.51 22.0 18.91 ;
    END
  END K<0>
END dotproduct_R

MACRO dotproduct_mid
  PIN GND
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 13.08 21.4 13.68 22.0 ;
    END
  END GND
  PIN out2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 17.05 21.4 17.65 22.0 ;
    END
  END out2
  PIN out1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 6.95 21.4 7.55 22.0 ;
    END
  END out1
  PIN phi2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 11.45 21.4 12.05 22.0 ;
    END
  END phi2
  PIN phi1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 2.1 21.4 2.7 22.0 ;
    END
  END phi1
  PIN Q<0>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 0.0 16.61 1.4 18.01 ;
    END
  END Q<0>
  PIN Q<3>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 0.0 4.01 1.4 5.41 ;
    END
  END Q<3>
  PIN Q<1>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 0.0 14.76 1.4 16.16 ;
    END
  END Q<1>
  PIN Q<2>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 0.0 5.86 1.4 7.26 ;
    END
  END Q<2>
  PIN K<2>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 20.6 9.31 22.0 10.71 ;
    END
  END K<2>
  PIN K<1>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 20.6 11.31 22.0 12.71 ;
    END
  END K<1>
  PIN K<3>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 20.6 0.56 22.0 1.96 ;
    END
  END K<3>
  PIN K<0>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 20.6 20.06 22.0 21.46 ;
    END
  END K<0>
END dotproduct_mid

MACRO dotproduct_L
  PIN K<0>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 20.6 20.05 22.0 21.45 ;
    END
  END K<0>
  PIN K<1>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 20.6 11.3 22.0 12.7 ;
    END
  END K<1>
  PIN Q<2>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 0.0 6.4 1.4 7.8 ;
    END
  END Q<2>
  PIN K<3>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 20.6 0.55 22.0 1.95 ;
    END
  END K<3>
  PIN Q<3>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 0.0 3.45 1.4 4.85 ;
    END
  END Q<3>
  PIN K<2>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 20.6 9.3 22.0 10.7 ;
    END
  END K<2>
  PIN Q<1>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 0.0 14.2 1.4 15.6 ;
    END
  END Q<1>
  PIN Q<0>
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
        RECT 0.0 17.15 1.4 18.55 ;
    END
  END Q<0>
  PIN GND
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 2.6 21.4 3.2 22.0 ;
    END
  END GND
  PIN phi1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 1.35 21.4 1.95 22.0 ;
    END
  END phi1
  PIN out2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 17.05 21.4 17.65 22.0 ;
    END
  END out2
  PIN phi2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 11.45 21.4 12.05 22.0 ;
    END
  END phi2
  PIN out1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 6.95 21.4 7.55 22.0 ;
    END
  END out1
END dotproduct_L

MACRO K_layer_output
  PIN GND
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 5.05 21.4 5.65 22.0 ;
    END
  END GND
END K_layer_output

END LIBRARY